`timescale 1ns / 1ns
module InstructionMemory(address,instruction);
  input[15:0] address;
  output[31:0]instruction;
  case address begin
endmodule
