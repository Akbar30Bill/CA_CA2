`timescale 1ns / 1ns
module Controller();
  
endmodule
